    package body package0 is
     function fn0 (param0 : bit_vector)
                       return bit is
      begin
        -- function code
      end fn0;
