entity HALFADD is
  port( a : in std_logic;
		b : in std_logic;
        sum : out std_logic;
        cary: out std_logic);
end HALFADD;
