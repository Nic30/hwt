package body package0 is
end package0;
